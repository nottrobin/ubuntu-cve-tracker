Candidate:
PublicDate:
References:
Description:
Ubuntu-Description:
Notes:
 leosilva> Issues that touch python_modules for spice in Xenial
 leosilva> need to be addressed in spice-protocol.
Bugs:
Priority: untriaged
Discovered-by:
Assigned-to:


Patches_spice-gtk:
upstream_spice-gtk: needs-triage
precise/esm_spice-gtk: DNE
trusty_spice-gtk: needs-triage
xenial_spice-gtk: needs-triage
bionic_spice-gtk: needs-triage
cosmic_spice-gtk: needs-triage
devel_spice-gtk: needs-triage

Patches_spice:
upstream_spice: needs-triage
precise/esm_spice: DNE
trusty_spice: needs-triage
xenial_spice: needs-triage
bionic_spice: needs-triage
cosmic_spice: needs-triage
devel_spice: needs-triage

Patches_spice-protocol:
upstream_spice-protocol: needs-triage
precise/esm_spice: DNE
trusty_spice-protocol: needs-triage
xenial_spice-protocol: needs-triage
bionic_spice-protocol: needs-triage
cosmic_spice-protocol: needs-triage
devel_spice-protocol: needs-triage
